library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity MemoryIO is

   PORT(
        -- Sistema
        CLK_SLOW : IN  STD_LOGIC;
        CLK_FAST : IN  STD_LOGIC;
        RST      : IN  STD_LOGIC;

        -- RAM 16K
        ADDRESS		: IN  STD_LOGIC_VECTOR (14 DOWNTO 0);
        INPUT		: IN  STD_LOGIC_VECTOR (15 DOWNTO 0);
        LOAD		: IN  STD_LOGIC ;
        OUTPUT		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);

        -- LCD EXTERNAL I/OS
        LCD_CS_N     : OUT   STD_LOGIC;
        LCD_D        : INOUT STD_LOGIC_VECTOR(15 downto 0);
        LCD_RD_N     : OUT   STD_LOGIC;
        LCD_RESET_N  : OUT   STD_LOGIC;
        LCD_RS       : OUT   STD_LOGIC;	-- (DCx) 0 : reg, 1: command
        LCD_WR_N     : OUT   STD_LOGIC;
        LCD_ON       : OUT   STD_LOGIC := '1';	-- liga e desliga o LCD
        LCD_INIT_OK  : OUT   STD_LOGIC;

        -- Switchs
        SW  : in std_logic_vector(9 downto 0);
        LED : OUT std_logic_vector(9 downto 0)

		);
end entity;


ARCHITECTURE logic OF MemoryIO IS

  component Screen is
      PORT(
          INPUT        : IN STD_LOGIC_VECTOR(15 downto 0);
          LOAD         : IN  STD_LOGIC;
          ADDRESS      : IN STD_LOGIC_VECTOR(13 downto 0);

          -- Sistema
          CLK_FAST : IN  STD_LOGIC;
          CLK_SLOW : IN  STD_LOGIC;
          RST 	   : IN  STD_LOGIC;

          -- LCD EXTERNAL I/OS
          LCD_INIT_OK  : OUT STD_LOGIC;
          LCD_CS_N     : OUT   STD_LOGIC;
          LCD_D        : INOUT STD_LOGIC_VECTOR(15 downto 0);
          LCD_RD_N     : OUT   STD_LOGIC;
          LCD_RESET_N  : OUT   STD_LOGIC;
          LCD_RS       : OUT   STD_LOGIC;	-- (DCx) 0 : reg, 1: command
          LCD_WR_N     : OUT   STD_LOGIC
          );
  end component;

  	component RAM16K IS
     	 PORT
      		(
          	address	: IN STD_LOGIC_VECTOR (13 DOWNTO 0);
          	clock		: IN STD_LOGIC  := '1';
          	data		: IN STD_LOGIC_VECTOR (15 DOWNTO 0);
         	wren		: IN STD_LOGIC ;
          	q		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
      		);
 	end component;

	component SCREEN IS
     	 PORT
      		(
          	address	: IN STD_LOGIC_VECTOR (13 DOWNTO 0);
          	clock_fast	: IN STD_LOGIC  := '1';
		clock_slow 	: IN STD_LOGIC  := '1';
          	load		: IN STD_LOGIC_VECTOR (15 DOWNTO 0);
         	input		: IN STD_LOGIC ;
          	LCD		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
      		);
 	end component;

  	component Register8 is
		port(

		clock:   in STD_LOGIC;
		input:   in STD_LOGIC_VECTOR(7 downto 0);
		load:    in STD_LOGIC;
		output: out  STD_LOGIC_VECTOR(7 downto 0)
		);
	end component;

BEGIN

m0: RAM16K port map (
	ADRESS => adress,
	CLK_FAST => clock,
	INPUT => data,
	LOAD => wren
   		     );
m1: SCREEN port map (
	ADRESS => adress,
	CLK_FAST => clock_fast,
	CLK_SLOW => clock_slow,
	LOAD => load,
	INPUT => input
		     );

m2: Register8 port map (
	CLK_FAST => clock,
	INPUT => input,
	LOAD => load,
		);

END logic;